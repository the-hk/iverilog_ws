// first_trial.v
module first_trial(
    input wire a,
    input wire b,
    output wire y
);

assign y = a 

endmodule
